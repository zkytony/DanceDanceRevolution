library verilog;
use verilog.vl_types.all;
entity score_counter_vlg_vec_tst is
end score_counter_vlg_vec_tst;
