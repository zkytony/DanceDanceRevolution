library verilog;
use verilog.vl_types.all;
entity score_keep_vlg_vec_tst is
end score_keep_vlg_vec_tst;
